
`timescale 1ns/1ns // set timescale
module fulladder(a,b,c,s, cout) ; // full adder circuit
input a , b, c ;  //declare inputs
output s, cout;  // declare outputs
 wire w1, w2, w3, w4;  // decalre wires
 xor #1     
 g1(w1, a, b), // xor a and b
 g2(s, w1, c);  // xor w1 and c
 and #1
 g3(w2, c, b), // c&b
 g4(w3, c, a), // c&a
 g5(w4, a, b); // a&b
 or #1
 g6(cout, w2, w3, w4); // w2|w3
 endmodule 
 
 module twotoonemux(a,b,s, f); // 2 to 1 mux circuit
 input a, b, s;  // declare inputs
 output f; // declare outputs
 wire w1, w2, w3;// declare wires
 not #1
 g1(w1, s); // ~s 
 and #1
 g2(w2, w1, a), // w1 & a
 g3(w3, s, b); // s&b
 or #1
 g4(f, w2, w3); // w2 | w3
 endmodule
 module fourtoonemux(a, b,c,d, s0, s1, f); // 4 to 1 mux circuit
 input a,b,c,d,s0,s1; // declare inputs
 output f; // declare outputs
wire w1,w2; // declare wires
twotoonemux m1(a,b,s1,w1); // uses 3 2 to 1 muxs using the output of the of the first 2 as inputs for the third mux
twotoonemux m2(c,d,s1,w2);
twotoonemux m3(w1,w2, s0,f);
endmodule
module bitalu(a,b,less,sub,cin,op0,op1, cout, out, set); // 1 bit alu circuit
input a,b,less,sub, cin, op0, op1; // decalre inputs
output cout, out, set; // declare outputs
wire w1, w2, w3, w4, w5, w6; // declare wires
and #1
g1(w1,a,b); // a&b
or #1
g2(w2,a,b); // a|b
not #1
g3(w3, b); //~b
twotoonemux m1(b,w3,sub,w4);    //two to one mux with b and w3 as inputs and sub as selector
fulladder f0(a,w4,cin,w5,cout); // full adder with a, w4, and cin as inputs
assign set = w5; // out of fulladder is set
fourtoonemux m2(w1,w2,w5,less,op0,op1, out); // 4 to 1 mux with w1, w2,w5, less as inputs and op0, op1 as selectors
endmodule

module alu(a,b,sub,op0,op1, out); //16 bit alu circuit
input [15:0] a,b;  // declare inputs
input op0,op1;
input sub;
output [15:0] out; //declare outputs
wire [16:0] w;// declare wires
wire se; // delcare set less wire
wire [14:0] c; // declare cin and cout wires
bitalu b1 (a[0],b[0],se,sub,sub,op0,op1,c[0], out[0], w[0]); // string together 16 1 bit alus with cout as cin for next alu, sub as cin for first and wire connecting the set of the last alu to the less of the first
bitalu b2(a[1],b[1],0,sub,c[0],op0,op1,c[1], out[1], w[1]);
bitalu b3(a[2],b[2],0,sub,c[1],op0,op1,c[2], out[2], w[2]);
bitalu b4(a[3],b[3],0,sub,c[2],op0,op1,c[3], out[3], w[3]);
bitalu b5(a[4],b[4],0,sub,c[3],op0,op1,c[4], out[4], w[4]);
bitalu b6(a[5],b[5],0,sub,c[4],op0,op1,c[5], out[5], w[5]);
bitalu b7(a[6],b[6],0,sub,c[5],op0,op1,c[6], out[6], w[6]);
bitalu b8(a[7],b[7],0,sub,c[6],op0,op1,c[7], out[7], w[7]);
bitalu b9(a[8],b[8],0,sub,c[7],op0,op1,c[8], out[8], w[8]);
bitalu b10(a[9],b[9],0,sub,c[8],op0,op1,c[9], out[9], w[9]);
bitalu b11(a[10],b[10],0,sub,c[9],op0,op1,c[10], out[10], w[10]);
bitalu b12(a[11],b[11],0,sub,c[10],op0,op1,c[11], out[11], w[11]);
bitalu b13(a[12],b[12],0,sub,c[11],op0,op1,c[12], out[12], w[12]);
bitalu b14(a[13],b[13],0,sub,c[12],op0,op1,c[13], out[13], w[13]);
bitalu b15(a[14],b[14],0,sub,c[13],op0,op1,c[14], out[14], w[14]);
bitalu b16(a[15],b[15],0,sub,c[14],op0,op1,w[15], out[15], se);
endmodule
module testbench(); //testbench creation
wire  [15:0] a,b;
wire sub , op0,op1;
wire [15:0] out;
testalu test(a,b,sub,op0,op1,out);  // connectinig alu to testbench alu
alu al(a,b,sub, op0, op1, out); 
endmodule

module testalu(a,b,sub,op0,op1,out); //outputs for testbench
output sub; // declare sub as output
input [15:0] out; // declare inputs
output [15:0] a,b; // declare outputs
output op0, op1;  // declare as output
reg op0, op1; //declare registers
reg [15:0] a,b;
reg sub;
initial
 begin
 $monitor($time, "a=%b, b=%b, sub=%b,op0=%b,op1=%b,out=%b",a,b,sub,op0,op1,out);
 $display($time, "a=%b, b=%b, sub=%b,op0=%b,op1=%b,out=%b",a,b,sub,op0,op1,out); 
#100 a=5053; b=1226; sub =0; op0=1; op1=0; // 5053 + 1226= 6279
#100 a=1844; b=2986; sub =0; op0=1; op1=0; // 1844 + 2986= 4830
#100 a=314; b=1930; sub =0; op0=0; op1=1; // 314 | 1930
#100 a=114; b=637; sub =1; op0=1; op1=0; // 114 - 637= -523
#100 a=149; b=7320; sub =1; op0=1; op1=1; // 149 < 7320
#100 a=5973; b=9361; sub =0; op0=0; op1=1; // 5973 | 9361
#100 a=4663; b=3853; sub =1; op0=1; op1=0; // 4663 - 3853= 810
#100 a=2088; b=346; sub =1; op0=1; op1=1; // 2088 < 346
#100 a=8067; b=2702; sub =1; op0=1; op1=0; // 8067 - 2702= 5365
#100 a=7209; b=8057; sub =0; op0=0; op1=0; // 7209 & 8057
#100 a=958; b=4924; sub =0; op0=1; op1=0; // 958 + 4924= 5882
#100 a=7834; b=8974; sub =1; op0=1; op1=1; // 7834 < 8974
#100 a=1470; b=6900; sub =1; op0=1; op1=0; // 1470 - 6900= -5430
#100 a=5658; b=7097; sub =0; op0=0; op1=1; // 5658 | 7097
#100 a=1633; b=9449; sub =1; op0=1; op1=1; // 1633 < 9449
#100 a=7364; b=4536; sub =1; op0=1; op1=0; // 7364 - 4536= 2828
#100 a=7520; b=4219; sub =0; op0=0; op1=1; // 7520 | 4219
#100 a=1465; b=900; sub =1; op0=1; op1=0; // 1465 - 900= 565
#100 a=7285; b=6024; sub =0; op0=0; op1=0; // 7285 & 6024
#100 a=9756; b=8784; sub =0; op0=1; op1=0; // 9756 + 8784= 18540
#100 a=7183; b=7899; sub =0; op0=0; op1=0; // 7183 & 7899
#100 a=7465; b=9175; sub =1; op0=1; op1=0; // 7465 - 9175= -1710
#100 a=5292; b=6468; sub =0; op0=0; op1=0; // 5292 & 6468
#100 a=4314; b=9641; sub =1; op0=1; op1=1; // 4314 < 9641
#100 a=5999; b=7799; sub =1; op0=1; op1=0; // 5999 - 7799= -1800
#100 a=5048; b=6262; sub =0; op0=1; op1=0; // 5048 + 6262= 11310
#100 a=4497; b=3592; sub =1; op0=1; op1=0; // 4497 - 3592= 905
#100 a=6705; b=8214; sub =0; op0=1; op1=0; // 6705 + 8214= 14919
#100 a=4140; b=2635; sub =0; op0=0; op1=0; // 4140 & 2635
#100 a=281; b=4518; sub =0; op0=0; op1=0; // 281 & 4518
#100 a=9390; b=8761; sub =1; op0=1; op1=0; // 9390 - 8761= 629
#100 a=3196; b=9677; sub =0; op0=0; op1=0; // 3196 & 9677
#100 a=6770; b=6444; sub =1; op0=1; op1=0; // 6770 - 6444= 326
#100 a=8623; b=6374; sub =1; op0=1; op1=1; // 8623 < 6374
#100 a=5144; b=9121; sub =0; op0=0; op1=0; // 5144 & 9121
#100 a=9349; b=2695; sub =0; op0=0; op1=0; // 9349 & 2695
#100 a=6212; b=379; sub =0; op0=1; op1=0; // 6212 + 379= 6591
#100 a=3465; b=9841; sub =1; op0=1; op1=0; // 3465 - 9841= -6376
#100 a=7931; b=8033; sub =1; op0=1; op1=0; // 7931 - 8033= -102
#100 a=4977; b=7712; sub =0; op0=0; op1=1; // 4977 | 7712
#100 a=20; b=5085; sub =1; op0=1; op1=0; // 20 - 5085= -5065
#100 a=7985; b=1101; sub =1; op0=1; op1=1; // 7985 < 1101
#100 a=739; b=6038; sub =0; op0=0; op1=0; // 739 & 6038
#100 a=4684; b=6247; sub =0; op0=0; op1=0; // 4684 & 6247
#100 a=7895; b=1495; sub =0; op0=0; op1=1; // 7895 | 1495
#100 a=455; b=9914; sub =1; op0=1; op1=1; // 455 < 9914
#100 a=395; b=9979; sub =0; op0=0; op1=1; // 395 | 9979
#100 a=3506; b=8460; sub =0; op0=0; op1=0; // 3506 & 8460
#100 a=3182; b=7065; sub =1; op0=1; op1=1; // 3182 < 7065
#100 a=3652; b=7259; sub =1; op0=1; op1=1; // 3652 < 7259
#100 a=3864; b=2435; sub =1; op0=1; op1=0; // 3864 - 2435= 1429
#100 a=4424; b=7302; sub =0; op0=1; op1=0; // 4424 + 7302= 11726
#100 a=7465; b=8699; sub =0; op0=0; op1=1; // 7465 | 8699
#100 a=4698; b=6375; sub =0; op0=0; op1=1; // 4698 | 6375
#100 a=7830; b=3607; sub =0; op0=0; op1=1; // 7830 | 3607
#100 a=4244; b=7035; sub =0; op0=1; op1=0; // 4244 + 7035= 11279
#100 a=1972; b=2981; sub =0; op0=1; op1=0; // 1972 + 2981= 4953
#100 a=6820; b=6787; sub =0; op0=0; op1=1; // 6820 | 6787
#100 a=2115; b=7454; sub =0; op0=0; op1=0; // 2115 & 7454
#100 a=3628; b=1184; sub =1; op0=1; op1=1; // 3628 < 1184
#100 a=6115; b=6382; sub =1; op0=1; op1=1; // 6115 < 6382
#100 a=8535; b=4278; sub =0; op0=0; op1=1; // 8535 | 4278
#100 a=8599; b=5848; sub =1; op0=1; op1=1; // 8599 < 5848
#100 a=7437; b=2496; sub =0; op0=1; op1=0; // 7437 + 2496= 9933
#100 a=1339; b=5972; sub =1; op0=1; op1=1; // 1339 < 5972
#100 a=1703; b=3134; sub =1; op0=1; op1=1; // 1703 < 3134
#100 a=1760; b=2018; sub =0; op0=0; op1=0; // 1760 & 2018
#100 a=2611; b=3627; sub =0; op0=0; op1=1; // 2611 | 3627
#100 a=44; b=9034; sub =0; op0=0; op1=0; // 44 & 9034
#100 a=1818; b=9469; sub =1; op0=1; op1=0; // 1818 - 9469= -7651
#100 a=52; b=3618; sub =1; op0=1; op1=0; // 52 - 3618= -3566
#100 a=4900; b=4451; sub =0; op0=0; op1=0; // 4900 & 4451
#100 a=1827; b=8134; sub =0; op0=0; op1=1; // 1827 | 8134
#100 a=1825; b=996; sub =0; op0=0; op1=0; // 1825 & 996
#100 a=5878; b=1737; sub =0; op0=1; op1=0; // 5878 + 1737= 7615
#100 a=3452; b=4224; sub =1; op0=1; op1=0; // 3452 - 4224= -772
#100 a=5512; b=7385; sub =0; op0=0; op1=0; // 5512 & 7385
#100 a=7490; b=7018; sub =0; op0=0; op1=0; // 7490 & 7018
#100 a=3260; b=3719; sub =0; op0=1; op1=0; // 3260 + 3719= 6979
#100 a=232; b=929; sub =0; op0=0; op1=1; // 232 | 929
#100 a=1722; b=8693; sub =0; op0=0; op1=0; // 1722 & 8693
#100 a=7486; b=7506; sub =1; op0=1; op1=0; // 7486 - 7506= -20
#100 a=4953; b=6442; sub =1; op0=1; op1=0; // 4953 - 6442= -1489
#100 a=4876; b=5725; sub =0; op0=1; op1=0; // 4876 + 5725= 10601
#100 a=1256; b=4402; sub =0; op0=1; op1=0; // 1256 + 4402= 5658
#100 a=8805; b=271; sub =0; op0=0; op1=1; // 8805 | 271
#100 a=4103; b=6931; sub =1; op0=1; op1=0; // 4103 - 6931= -2828
#100 a=5314; b=142; sub =1; op0=1; op1=0; // 5314 - 142= 5172
#100 a=425; b=7197; sub =0; op0=0; op1=0; // 425 & 7197
#100 a=2202; b=4233; sub =0; op0=0; op1=0; // 2202 & 4233
#100 a=5799; b=5525; sub =1; op0=1; op1=0; // 5799 - 5525= 274
#100 a=865; b=7351; sub =1; op0=1; op1=1; // 865 < 7351
#100 a=396; b=5711; sub =1; op0=1; op1=0; // 396 - 5711= -5315
#100 a=3116; b=1616; sub =0; op0=0; op1=1; // 3116 | 1616
#100 a=1419; b=1567; sub =0; op0=0; op1=0; // 1419 & 1567
#100 a=9213; b=5984; sub =1; op0=1; op1=1; // 9213 < 5984
#100 a=3936; b=522; sub =0; op0=0; op1=0; // 3936 & 522
#100 a=1541; b=3993; sub =0; op0=0; op1=1; // 1541 | 3993
#100 a=6181; b=2585; sub =0; op0=0; op1=1; // 6181 | 2585
#100 a=3349; b=8278; sub =1; op0=1; op1=1; // 3349 < 8278
#100 a=7870; b=9555; sub =0; op0=0; op1=0; // 7870 & 9555
#100 a=3155; b=365; sub =0; op0=0; op1=0; // 3155 & 365
#100 a=6077; b=5148; sub =1; op0=1; op1=0; // 6077 - 5148= 929
#100 a=6531; b=3779; sub =1; op0=1; op1=1; // 6531 < 3779
#100 a=4210; b=2371; sub =0; op0=0; op1=1; // 4210 | 2371
#100 a=4069; b=7793; sub =1; op0=1; op1=0; // 4069 - 7793= -3724
#100 a=4964; b=811; sub =0; op0=0; op1=1; // 4964 | 811
#100 a=175; b=4648; sub =1; op0=1; op1=0; // 175 - 4648= -4473
#100 a=1127; b=4361; sub =1; op0=1; op1=0; // 1127 - 4361= -3234
#100 a=6528; b=2523; sub =1; op0=1; op1=0; // 6528 - 2523= 4005
#100 a=163; b=9680; sub =0; op0=1; op1=0; // 163 + 9680= 9843
#100 a=1727; b=5180; sub =1; op0=1; op1=0; // 1727 - 5180= -3453
#100 a=166; b=9819; sub =0; op0=1; op1=0; // 166 + 9819= 9985
#100 a=5184; b=6407; sub =0; op0=0; op1=1; // 5184 | 6407
#100 a=3734; b=4622; sub =0; op0=1; op1=0; // 3734 + 4622= 8356
#100 a=9730; b=9766; sub =0; op0=0; op1=1; // 9730 | 9766
#100 a=5780; b=1925; sub =0; op0=0; op1=1; // 5780 | 1925
#100 a=5264; b=3318; sub =1; op0=1; op1=0; // 5264 - 3318= 1946
#100 a=6688; b=3436; sub =0; op0=1; op1=0; // 6688 + 3436= 10124
#100 a=6408; b=7861; sub =1; op0=1; op1=1; // 6408 < 7861
#100 a=5297; b=3305; sub =1; op0=1; op1=1; // 5297 < 3305
#100 a=8363; b=7267; sub =1; op0=1; op1=0; // 8363 - 7267= 1096
#100 a=3377; b=1029; sub =1; op0=1; op1=0; // 3377 - 1029= 2348
#100 a=6886; b=3521; sub =1; op0=1; op1=0; // 6886 - 3521= 3365
#100 a=1646; b=7489; sub =1; op0=1; op1=0; // 1646 - 7489= -5843
#100 a=5816; b=7998; sub =1; op0=1; op1=0; // 5816 - 7998= -2182
#100 a=9866; b=1012; sub =0; op0=1; op1=0; // 9866 + 1012= 10878
#100 a=6342; b=6574; sub =0; op0=0; op1=0; // 6342 & 6574
#100 a=1294; b=7822; sub =1; op0=1; op1=1; // 1294 < 7822
#100 a=5584; b=3500; sub =1; op0=1; op1=0; // 5584 - 3500= 2084
#100 a=8586; b=4617; sub =0; op0=0; op1=0; // 8586 & 4617
#100 a=4236; b=4378; sub =0; op0=1; op1=0; // 4236 + 4378= 8614
#100 a=9966; b=7317; sub =0; op0=0; op1=1; // 9966 | 7317
#100 a=578; b=8819; sub =0; op0=0; op1=0; // 578 & 8819
#100 a=9266; b=6329; sub =1; op0=1; op1=1; // 9266 < 6329
#100 a=1491; b=1910; sub =0; op0=0; op1=0; // 1491 & 1910
#100 a=3465; b=7928; sub =1; op0=1; op1=0; // 3465 - 7928= -4463
#100 a=7631; b=1766; sub =1; op0=1; op1=1; // 7631 < 1766
#100 a=9; b=4474; sub =0; op0=0; op1=1; // 9 | 4474
#100 a=2612; b=8311; sub =1; op0=1; op1=1; // 2612 < 8311
#100 a=7283; b=3953; sub =0; op0=0; op1=0; // 7283 & 3953
#100 a=5935; b=430; sub =0; op0=0; op1=1; // 5935 | 430
#100 a=1308; b=3912; sub =0; op0=1; op1=0; // 1308 + 3912= 5220
#100 a=1802; b=5900; sub =1; op0=1; op1=1; // 1802 < 5900
#100 a=417; b=2296; sub =0; op0=0; op1=0; // 417 & 2296
#100 a=7103; b=1364; sub =0; op0=0; op1=1; // 7103 | 1364
#100 a=2742; b=2188; sub =0; op0=1; op1=0; // 2742 + 2188= 4930
#100 a=1391; b=1637; sub =1; op0=1; op1=0; // 1391 - 1637= -246
#100 a=7738; b=9061; sub =0; op0=1; op1=0; // 7738 + 9061= 16799
#100 a=6142; b=6756; sub =0; op0=0; op1=0; // 6142 & 6756
#100 a=4799; b=4568; sub =0; op0=0; op1=1; // 4799 | 4568
#100 a=263; b=4132; sub =0; op0=1; op1=0; // 263 + 4132= 4395
#100 a=197; b=9607; sub =0; op0=1; op1=0; // 197 + 9607= 9804
#100 a=5100; b=1700; sub =0; op0=0; op1=0; // 5100 & 1700
#100 a=2389; b=657; sub =0; op0=0; op1=0; // 2389 & 657
#100 a=8020; b=2930; sub =0; op0=1; op1=0; // 8020 + 2930= 10950
#100 a=9354; b=7344; sub =0; op0=1; op1=0; // 9354 + 7344= 16698
#100 a=3916; b=9919; sub =1; op0=1; op1=0; // 3916 - 9919= -6003
#100 a=4046; b=5828; sub =0; op0=0; op1=1; // 4046 | 5828
#100 a=3456; b=1536; sub =1; op0=1; op1=0; // 3456 - 1536= 1920
#100 a=1966; b=8858; sub =1; op0=1; op1=0; // 1966 - 8858= -6892
#100 a=5070; b=2010; sub =0; op0=1; op1=0; // 5070 + 2010= 7080
#100 a=5905; b=7639; sub =0; op0=1; op1=0; // 5905 + 7639= 13544
#100 a=4567; b=2928; sub =1; op0=1; op1=0; // 4567 - 2928= 1639
#100 a=8977; b=1437; sub =1; op0=1; op1=0; // 8977 - 1437= 7540
#100 a=4909; b=2342; sub =0; op0=0; op1=1; // 4909 | 2342
#100 a=8148; b=3564; sub =0; op0=0; op1=1; // 8148 | 3564
#100 a=5609; b=9399; sub =1; op0=1; op1=0; // 5609 - 9399= -3790
#100 a=2561; b=494; sub =0; op0=1; op1=0; // 2561 + 494= 3055
#100 a=7919; b=7381; sub =1; op0=1; op1=0; // 7919 - 7381= 538
#100 a=3646; b=410; sub =0; op0=0; op1=1; // 3646 | 410
#100 a=9275; b=9471; sub =0; op0=0; op1=0; // 9275 & 9471
#100 a=1196; b=1978; sub =1; op0=1; op1=1; // 1196 < 1978
#100 a=7402; b=9893; sub =0; op0=0; op1=0; // 7402 & 9893
#100 a=3826; b=1530; sub =0; op0=0; op1=0; // 3826 & 1530
#100 a=7978; b=6610; sub =0; op0=1; op1=0; // 7978 + 6610= 14588
#100 a=5964; b=8707; sub =0; op0=0; op1=1; // 5964 | 8707
#100 a=3431; b=796; sub =0; op0=1; op1=0; // 3431 + 796= 4227
#100 a=1990; b=4065; sub =0; op0=0; op1=0; // 1990 & 4065
#100 a=1638; b=7444; sub =0; op0=0; op1=0; // 1638 & 7444
#100 a=2738; b=9971; sub =0; op0=1; op1=0; // 2738 + 9971= 12709
#100 a=1243; b=8594; sub =1; op0=1; op1=1; // 1243 < 8594
#100 a=2341; b=4858; sub =1; op0=1; op1=0; // 2341 - 4858= -2517
#100 a=7953; b=1169; sub =0; op0=0; op1=0; // 7953 & 1169
#100 a=6651; b=1780; sub =0; op0=0; op1=1; // 6651 | 1780
#100 a=4169; b=3021; sub =1; op0=1; op1=0; // 4169 - 3021= 1148
#100 a=2939; b=6292; sub =0; op0=0; op1=0; // 2939 & 6292
#100 a=9470; b=9445; sub =1; op0=1; op1=1; // 9470 < 9445
#100 a=9745; b=4459; sub =1; op0=1; op1=1; // 9745 < 4459
#100 a=6725; b=6869; sub =1; op0=1; op1=0; // 6725 - 6869= -144
#100 a=4667; b=1079; sub =1; op0=1; op1=1; // 4667 < 1079
#100 a=8270; b=8625; sub =1; op0=1; op1=0; // 8270 - 8625= -355
#100 a=5487; b=1428; sub =0; op0=0; op1=0; // 5487 & 1428
#100 a=6326; b=7977; sub =0; op0=0; op1=1; // 6326 | 7977
#100 a=5399; b=9220; sub =0; op0=0; op1=1; // 5399 | 9220
#100 a=1328; b=6013; sub =1; op0=1; op1=1; // 1328 < 6013
#100 a=6410; b=4138; sub =0; op0=1; op1=0; // 6410 + 4138= 10548
#100 a=1823; b=1281; sub =1; op0=1; op1=1; // 1823 < 1281
#100 a=7024; b=7066; sub =1; op0=1; op1=0; // 7024 - 7066= -42
#100 a=7840; b=3297; sub =1; op0=1; op1=0; // 7840 - 3297= 4543
#100 a=7070; b=3012; sub =0; op0=0; op1=1; // 7070 | 3012
#100 a=6367; b=8367; sub =1; op0=1; op1=0; // 6367 - 8367= -2000
#100 a=3227; b=5738; sub =1; op0=1; op1=0; // 3227 - 5738= -2511
#100 a=5645; b=3924; sub =0; op0=0; op1=0; // 5645 & 3924
#100 a=8422; b=4382; sub =1; op0=1; op1=1; // 8422 < 4382
#100 a=2636; b=7601; sub =1; op0=1; op1=0; // 2636 - 7601= -4965
#100 a=639; b=4599; sub =1; op0=1; op1=1; // 639 < 4599
#100 a=4082; b=8421; sub =0; op0=0; op1=0; // 4082 & 8421
#100 a=8003; b=9026; sub =0; op0=0; op1=1; // 8003 | 9026
#100 a=6801; b=3455; sub =1; op0=1; op1=0; // 6801 - 3455= 3346
#100 a=2882; b=4412; sub =1; op0=1; op1=1; // 2882 < 4412
#100 a=6922; b=1463; sub =1; op0=1; op1=0; // 6922 - 1463= 5459
#100 a=4413; b=3604; sub =1; op0=1; op1=0; // 4413 - 3604= 809
#100 a=535; b=9728; sub =0; op0=0; op1=0; // 535 & 9728
#100 a=4002; b=9886; sub =1; op0=1; op1=0; // 4002 - 9886= -5884
#100 a=9299; b=9939; sub =1; op0=1; op1=0; // 9299 - 9939= -640
#100 a=7938; b=2844; sub =0; op0=1; op1=0; // 7938 + 2844= 10782
#100 a=6090; b=6472; sub =0; op0=0; op1=1; // 6090 | 6472
#100 a=8732; b=8609; sub =0; op0=0; op1=0; // 8732 & 8609
#100 a=6567; b=1272; sub =0; op0=0; op1=0; // 6567 & 1272
#100 a=7457; b=3390; sub =0; op0=1; op1=0; // 7457 + 3390= 10847
#100 a=5160; b=3361; sub =1; op0=1; op1=0; // 5160 - 3361= 1799
#100 a=1513; b=2870; sub =1; op0=1; op1=1; // 1513 < 2870
#100 a=9901; b=8255; sub =0; op0=1; op1=0; // 9901 + 8255= 18156
#100 a=4807; b=8665; sub =1; op0=1; op1=0; // 4807 - 8665= -3858
#100 a=6985; b=4605; sub =0; op0=0; op1=0; // 6985 & 4605
#100 a=4968; b=9890; sub =1; op0=1; op1=1; // 4968 < 9890
#100 a=431; b=9003; sub =0; op0=0; op1=0; // 431 & 9003
#100 a=3824; b=897; sub =0; op0=0; op1=0; // 3824 & 897
#100 a=7428; b=6180; sub =1; op0=1; op1=1; // 7428 < 6180
#100 a=6080; b=5752; sub =1; op0=1; op1=0; // 6080 - 5752= 328
#100 a=4071; b=6086; sub =1; op0=1; op1=1; // 4071 < 6086
#100 a=324; b=1410; sub =1; op0=1; op1=1; // 324 < 1410
#100 a=9460; b=9153; sub =1; op0=1; op1=1; // 9460 < 9153
#100 a=79; b=580; sub =1; op0=1; op1=1; // 79 < 580
#100 a=1420; b=8704; sub =0; op0=0; op1=0; // 1420 & 8704
#100 a=2941; b=1154; sub =1; op0=1; op1=1; // 2941 < 1154
#100 a=4924; b=3601; sub =0; op0=0; op1=0; // 4924 & 3601
#100 a=4087; b=4302; sub =0; op0=0; op1=1; // 4087 | 4302
#100 a=8304; b=5891; sub =1; op0=1; op1=0; // 8304 - 5891= 2413
#100 a=7786; b=1435; sub =1; op0=1; op1=1; // 7786 < 1435
#100 a=600; b=8522; sub =0; op0=1; op1=0; // 600 + 8522= 9122
#100 a=9960; b=6710; sub =1; op0=1; op1=0; // 9960 - 6710= 3250
#100 a=8556; b=7380; sub =1; op0=1; op1=1; // 8556 < 7380
#100 a=1626; b=1908; sub =0; op0=1; op1=0; // 1626 + 1908= 3534
#100 a=2209; b=7299; sub =1; op0=1; op1=0; // 2209 - 7299= -5090
#100 a=9570; b=9900; sub =1; op0=1; op1=0; // 9570 - 9900= -330
#100 a=4022; b=9863; sub =0; op0=0; op1=0; // 4022 & 9863
#100 a=4338; b=4506; sub =0; op0=0; op1=1; // 4338 | 4506
#100 a=5298; b=6230; sub =1; op0=1; op1=1; // 5298 < 6230
#100 a=652; b=7453; sub =0; op0=1; op1=0; // 652 + 7453= 8105
#100 a=8281; b=5271; sub =0; op0=0; op1=1; // 8281 | 5271
#100 a=4464; b=1489; sub =0; op0=0; op1=1; // 4464 | 1489
#100 a=9404; b=9580; sub =1; op0=1; op1=1; // 9404 < 9580
#100 a=4260; b=4177; sub =1; op0=1; op1=0; // 4260 - 4177= 83
#100 a=6994; b=8303; sub =1; op0=1; op1=0; // 6994 - 8303= -1309
#100 a=7091; b=642; sub =0; op0=0; op1=0; // 7091 & 642
#100 a=5484; b=2389; sub =0; op0=0; op1=0; // 5484 & 2389
#100 a=8382; b=3370; sub =0; op0=0; op1=0; // 8382 & 3370
#100 a=1813; b=2018; sub =1; op0=1; op1=0; // 1813 - 2018= -205
#100 a=3; b=5590; sub =0; op0=1; op1=0; // 3 + 5590= 5593
#100 a=4088; b=8456; sub =1; op0=1; op1=1; // 4088 < 8456
#100 a=2336; b=5266; sub =0; op0=0; op1=0; // 2336 & 5266
#100 a=6834; b=7293; sub =1; op0=1; op1=1; // 6834 < 7293
#100 a=4474; b=41; sub =0; op0=1; op1=0; // 4474 + 41= 4515
#100 a=2629; b=125; sub =0; op0=0; op1=1; // 2629 | 125
#100 a=96; b=2741; sub =0; op0=0; op1=1; // 96 | 2741
#100 a=9721; b=7495; sub =1; op0=1; op1=0; // 9721 - 7495= 2226
#100 a=6347; b=8576; sub =1; op0=1; op1=1; // 6347 < 8576
#100 a=7221; b=5666; sub =1; op0=1; op1=0; // 7221 - 5666= 1555
#100 a=5090; b=6867; sub =1; op0=1; op1=1; // 5090 < 6867
#100 a=9481; b=9214; sub =0; op0=0; op1=1; // 9481 | 9214
#100 a=2602; b=6128; sub =1; op0=1; op1=0; // 2602 - 6128= -3526
#100 a=8644; b=7243; sub =1; op0=1; op1=0; // 8644 - 7243= 1401
#100 a=9623; b=6166; sub =1; op0=1; op1=1; // 9623 < 6166
#100 a=1804; b=1207; sub =1; op0=1; op1=0; // 1804 - 1207= 597
#100 a=7109; b=1499; sub =1; op0=1; op1=1; // 7109 < 1499
#100 a=5758; b=8941; sub =0; op0=1; op1=0; // 5758 + 8941= 14699
#100 a=5063; b=248; sub =0; op0=0; op1=1; // 5063 | 248
#100 a=6224; b=8866; sub =0; op0=1; op1=0; // 6224 + 8866= 15090
#100 a=6625; b=3405; sub =1; op0=1; op1=0; // 6625 - 3405= 3220
#100 a=5586; b=8221; sub =0; op0=0; op1=1; // 5586 | 8221
#100 a=84; b=1011; sub =0; op0=0; op1=0; // 84 & 1011
#100 a=4680; b=8943; sub =1; op0=1; op1=0; // 4680 - 8943= -4263
#100 a=2657; b=1448; sub =1; op0=1; op1=0; // 2657 - 1448= 1209
#100 a=6240; b=7490; sub =0; op0=0; op1=0; // 6240 & 7490
#100 a=2007; b=4033; sub =1; op0=1; op1=0; // 2007 - 4033= -2026
#100 a=9188; b=6452; sub =0; op0=0; op1=1; // 9188 | 6452
#100 a=4930; b=1358; sub =0; op0=0; op1=1; // 4930 | 1358
#100 a=3650; b=6422; sub =0; op0=1; op1=0; // 3650 + 6422= 10072
#100 a=4383; b=8978; sub =1; op0=1; op1=1; // 4383 < 8978
#100 a=2581; b=6354; sub =1; op0=1; op1=1; // 2581 < 6354
#100 a=1027; b=3522; sub =0; op0=1; op1=0; // 1027 + 3522= 4549
#100 a=8125; b=5006; sub =1; op0=1; op1=1; // 8125 < 5006
#100 a=3572; b=4975; sub =0; op0=0; op1=1; // 3572 | 4975
#100 a=6428; b=3192; sub =0; op0=0; op1=1; // 6428 | 3192
#100 a=5458; b=9270; sub =0; op0=0; op1=0; // 5458 & 9270
#100 a=3628; b=9550; sub =1; op0=1; op1=0; // 3628 - 9550= -5922
#100 a=6242; b=6481; sub =1; op0=1; op1=1; // 6242 < 6481
#100 a=4701; b=6194; sub =0; op0=0; op1=1; // 4701 | 6194
#100 a=3266; b=7127; sub =0; op0=0; op1=1; // 3266 | 7127
#100 a=6454; b=8447; sub =1; op0=1; op1=1; // 6454 < 8447
#100 a=360; b=9683; sub =0; op0=0; op1=1; // 360 | 9683
#100 a=5809; b=5057; sub =1; op0=1; op1=0; // 5809 - 5057= 752
#100 a=5451; b=7679; sub =0; op0=1; op1=0; // 5451 + 7679= 13130
#100 a=8888; b=2987; sub =1; op0=1; op1=1; // 8888 < 2987
#100 a=2945; b=8610; sub =0; op0=0; op1=1; // 2945 | 8610
#100 a=8464; b=1903; sub =1; op0=1; op1=1; // 8464 < 1903
#100 a=5821; b=4530; sub =0; op0=0; op1=0; // 5821 & 4530
#100 a=331; b=9801; sub =1; op0=1; op1=1; // 331 < 9801
#100 a=1101; b=2517; sub =1; op0=1; op1=0; // 1101 - 2517= -1416
#100 a=8682; b=3998; sub =0; op0=1; op1=0; // 8682 + 3998= 12680
#100 a=9768; b=4027; sub =1; op0=1; op1=0; // 9768 - 4027= 5741
#100 a=3574; b=5616; sub =1; op0=1; op1=1; // 3574 < 5616
#100 a=7062; b=7063; sub =0; op0=1; op1=0; // 7062 + 7063= 14125
#100 a=3457; b=5811; sub =0; op0=0; op1=0; // 3457 & 5811
#100 a=4462; b=1605; sub =0; op0=1; op1=0; // 4462 + 1605= 6067
#100 a=7956; b=2071; sub =0; op0=0; op1=1; // 7956 | 2071
#100 a=3029; b=9177; sub =0; op0=0; op1=1; // 3029 | 9177
#100 a=9490; b=4167; sub =0; op0=0; op1=0; // 9490 & 4167
#100 a=7957; b=2037; sub =0; op0=0; op1=1; // 7957 | 2037
#100 a=1263; b=9718; sub =1; op0=1; op1=0; // 1263 - 9718= -8455
#100 a=245; b=3532; sub =0; op0=1; op1=0; // 245 + 3532= 3777
#100 a=2238; b=8768; sub =0; op0=0; op1=1; // 2238 | 8768
#100 a=2399; b=2535; sub =0; op0=0; op1=0; // 2399 & 2535
#100 a=5451; b=3057; sub =0; op0=1; op1=0; // 5451 + 3057= 8508
#100 a=7235; b=5771; sub =0; op0=0; op1=0; // 7235 & 5771
#100 a=6798; b=3306; sub =1; op0=1; op1=1; // 6798 < 3306
#100 a=3120; b=9934; sub =0; op0=0; op1=0; // 3120 & 9934
#100 a=1191; b=9004; sub =1; op0=1; op1=1; // 1191 < 9004
#100 a=3543; b=783; sub =1; op0=1; op1=0; // 3543 - 783= 2760
#100 a=7709; b=5370; sub =0; op0=0; op1=0; // 7709 & 5370
#100 a=5809; b=7326; sub =1; op0=1; op1=1; // 5809 < 7326
#100 a=6442; b=680; sub =0; op0=0; op1=0; // 6442 & 680
#100 a=5420; b=9760; sub =1; op0=1; op1=1; // 5420 < 9760
#100 a=1410; b=726; sub =0; op0=1; op1=0; // 1410 + 726= 2136
#100 a=1638; b=4726; sub =1; op0=1; op1=0; // 1638 - 4726= -3088
#100 a=1280; b=7467; sub =1; op0=1; op1=1; // 1280 < 7467
#100 a=9916; b=5435; sub =0; op0=0; op1=0; // 9916 & 5435
#100 a=4831; b=2805; sub =0; op0=0; op1=1; // 4831 | 2805
#100 a=8066; b=3457; sub =1; op0=1; op1=1; // 8066 < 3457
#100 a=4134; b=1822; sub =0; op0=0; op1=0; // 4134 & 1822
#100 a=213; b=5985; sub =0; op0=0; op1=1; // 213 | 5985
#100 a=4491; b=8531; sub =1; op0=1; op1=0; // 4491 - 8531= -4040
#100 a=9390; b=8356; sub =0; op0=1; op1=0; // 9390 + 8356= 17746
#100 a=7477; b=8619; sub =1; op0=1; op1=0; // 7477 - 8619= -1142
#100 a=2670; b=7048; sub =0; op0=1; op1=0; // 2670 + 7048= 9718
#100 a=3598; b=9075; sub =1; op0=1; op1=0; // 3598 - 9075= -5477
#100 a=9272; b=883; sub =1; op0=1; op1=1; // 9272 < 883
#100 a=7903; b=6680; sub =0; op0=1; op1=0; // 7903 + 6680= 14583
#100 a=4802; b=2987; sub =1; op0=1; op1=0; // 4802 - 2987= 1815
#100 a=7998; b=998; sub =0; op0=0; op1=0; // 7998 & 998
#100 a=7899; b=5758; sub =1; op0=1; op1=0; // 7899 - 5758= 2141
#100 a=7025; b=6449; sub =1; op0=1; op1=0; // 7025 - 6449= 576
#100 a=2012; b=9894; sub =0; op0=0; op1=1; // 2012 | 9894
#100 a=4618; b=9644; sub =1; op0=1; op1=1; // 4618 < 9644
#100 a=5078; b=3033; sub =0; op0=0; op1=0; // 5078 & 3033
#100 a=3300; b=8451; sub =1; op0=1; op1=0; // 3300 - 8451= -5151
#100 a=4226; b=8889; sub =1; op0=1; op1=0; // 4226 - 8889= -4663
#100 a=6879; b=7193; sub =0; op0=0; op1=1; // 6879 | 7193
#100 a=1377; b=2435; sub =1; op0=1; op1=0; // 1377 - 2435= -1058
#100 a=8567; b=5647; sub =0; op0=0; op1=0; // 8567 & 5647
#100 a=659; b=6159; sub =0; op0=1; op1=0; // 659 + 6159= 6818
#100 a=182; b=1890; sub =0; op0=0; op1=0; // 182 & 1890
#100 a=2843; b=1108; sub =0; op0=1; op1=0; // 2843 + 1108= 3951
#100 a=7072; b=9436; sub =1; op0=1; op1=1; // 7072 < 9436
#100 a=5085; b=3786; sub =0; op0=0; op1=1; // 5085 | 3786
#100 a=5426; b=6642; sub =0; op0=0; op1=1; // 5426 | 6642
#100 a=8242; b=8894; sub =0; op0=1; op1=0; // 8242 + 8894= 17136
#100 a=481; b=8925; sub =0; op0=0; op1=0; // 481 & 8925
#100 a=1583; b=6333; sub =0; op0=0; op1=0; // 1583 & 6333
#100 a=8907; b=4040; sub =1; op0=1; op1=1; // 8907 < 4040
#100 a=6102; b=8851; sub =0; op0=1; op1=0; // 6102 + 8851= 14953
#100 a=9090; b=3220; sub =0; op0=0; op1=0; // 9090 & 3220
#100 a=4340; b=227; sub =1; op0=1; op1=1; // 4340 < 227
#100 a=9169; b=4552; sub =0; op0=1; op1=0; // 9169 + 4552= 13721
#100 a=3780; b=7860; sub =0; op0=0; op1=0; // 3780 & 7860
#100 a=6085; b=9329; sub =0; op0=1; op1=0; // 6085 + 9329= 15414
#100 a=8488; b=7255; sub =1; op0=1; op1=1; // 8488 < 7255
#100 a=1083; b=5916; sub =0; op0=0; op1=0; // 1083 & 5916
#100 a=8046; b=5692; sub =1; op0=1; op1=1; // 8046 < 5692
#100 a=2853; b=3054; sub =0; op0=1; op1=0; // 2853 + 3054= 5907
#100 a=8774; b=590; sub =0; op0=1; op1=0; // 8774 + 590= 9364
#100 a=1563; b=8012; sub =0; op0=0; op1=1; // 1563 | 8012
#100 a=9524; b=5937; sub =1; op0=1; op1=0; // 9524 - 5937= 3587
#100 a=2761; b=3734; sub =0; op0=0; op1=1; // 2761 | 3734
#100 a=5567; b=9680; sub =0; op0=1; op1=0; // 5567 + 9680= 15247
#100 a=8593; b=547; sub =0; op0=0; op1=0; // 8593 & 547
#100 a=9722; b=9788; sub =1; op0=1; op1=0; // 9722 - 9788= -66
#100 a=132; b=2339; sub =1; op0=1; op1=1; // 132 < 2339
#100 a=6542; b=2989; sub =0; op0=1; op1=0; // 6542 + 2989= 9531
#100 a=9542; b=8240; sub =1; op0=1; op1=1; // 9542 < 8240
#100 a=3770; b=2201; sub =0; op0=1; op1=0; // 3770 + 2201= 5971
#100 a=9999; b=697; sub =0; op0=1; op1=0; // 9999 + 697= 10696
#100 a=3941; b=8652; sub =1; op0=1; op1=1; // 3941 < 8652
#100 a=8178; b=7393; sub =0; op0=0; op1=0; // 8178 & 7393
#100 a=6520; b=1434; sub =0; op0=0; op1=1; // 6520 | 1434
#100 a=3814; b=3726; sub =0; op0=0; op1=0; // 3814 & 3726
#100 a=7619; b=4365; sub =0; op0=0; op1=0; // 7619 & 4365
#100 a=2327; b=5294; sub =1; op0=1; op1=1; // 2327 < 5294
#100 a=4107; b=1639; sub =1; op0=1; op1=1; // 4107 < 1639
#100 a=3695; b=1482; sub =1; op0=1; op1=0; // 3695 - 1482= 2213
#100 a=6886; b=9499; sub =1; op0=1; op1=1; // 6886 < 9499
#100 a=3214; b=9835; sub =1; op0=1; op1=0; // 3214 - 9835= -6621
#100 a=936; b=8372; sub =0; op0=0; op1=1; // 936 | 8372
#100 a=9301; b=7381; sub =0; op0=0; op1=1; // 9301 | 7381
#100 a=8212; b=4887; sub =0; op0=0; op1=1; // 8212 | 4887
#100 a=3862; b=4184; sub =1; op0=1; op1=1; // 3862 < 4184
#100 a=2846; b=328; sub =1; op0=1; op1=0; // 2846 - 328= 2518
#100 a=5887; b=6497; sub =0; op0=0; op1=0; // 5887 & 6497
#100 a=537; b=6381; sub =0; op0=0; op1=0; // 537 & 6381
#100 a=5237; b=2686; sub =0; op0=0; op1=1; // 5237 | 2686
#100 a=5931; b=9866; sub =0; op0=0; op1=1; // 5931 | 9866
#100 a=1882; b=190; sub =1; op0=1; op1=1; // 1882 < 190
#100 a=9818; b=8981; sub =1; op0=1; op1=0; // 9818 - 8981= 837
#100 a=9651; b=2181; sub =1; op0=1; op1=1; // 9651 < 2181
#100 a=9618; b=6117; sub =0; op0=1; op1=0; // 9618 + 6117= 15735
#100 a=2598; b=7541; sub =0; op0=0; op1=0; // 2598 & 7541
#100 a=2012; b=4182; sub =1; op0=1; op1=0; // 2012 - 4182= -2170
#100 a=8723; b=7680; sub =0; op0=0; op1=1; // 8723 | 7680
#100 a=123; b=5905; sub =0; op0=0; op1=1; // 123 | 5905
#100 a=2264; b=2813; sub =1; op0=1; op1=0; // 2264 - 2813= -549
#100 a=9227; b=74; sub =0; op0=0; op1=0; // 9227 & 74
#100 a=7032; b=3802; sub =0; op0=1; op1=0; // 7032 + 3802= 10834
#100 a=5397; b=8294; sub =1; op0=1; op1=1; // 5397 < 8294
#100 a=1622; b=8430; sub =1; op0=1; op1=1; // 1622 < 8430
#100 a=1222; b=5233; sub =0; op0=0; op1=1; // 1222 | 5233
#100 a=2752; b=7172; sub =0; op0=0; op1=1; // 2752 | 7172
#100 a=6502; b=5671; sub =0; op0=0; op1=1; // 6502 | 5671
#100 a=8447; b=5401; sub =0; op0=0; op1=0; // 8447 & 5401
#100 a=706; b=128; sub =0; op0=0; op1=0; // 706 & 128
#100 a=9630; b=9211; sub =1; op0=1; op1=0; // 9630 - 9211= 419
#100 a=666; b=7934; sub =0; op0=1; op1=0; // 666 + 7934= 8600
#100 a=1151; b=1701; sub =0; op0=0; op1=1; // 1151 | 1701
#100 a=8081; b=2464; sub =1; op0=1; op1=0; // 8081 - 2464= 5617
#100 a=9228; b=8567; sub =0; op0=0; op1=0; // 9228 & 8567
#100 a=4666; b=6937; sub =0; op0=0; op1=1; // 4666 | 6937
#100 a=8719; b=2330; sub =1; op0=1; op1=0; // 8719 - 2330= 6389
#100 a=7647; b=6469; sub =1; op0=1; op1=0; // 7647 - 6469= 1178
#100 a=6403; b=7768; sub =0; op0=1; op1=0; // 6403 + 7768= 14171
#100 a=1507; b=1725; sub =1; op0=1; op1=0; // 1507 - 1725= -218
#100 a=5856; b=7135; sub =0; op0=0; op1=0; // 5856 & 7135
#100 a=7683; b=8921; sub =0; op0=0; op1=1; // 7683 | 8921
#100 a=4827; b=6572; sub =1; op0=1; op1=0; // 4827 - 6572= -1745
#100 a=1740; b=5688; sub =1; op0=1; op1=1; // 1740 < 5688
#100 a=8979; b=6709; sub =1; op0=1; op1=0; // 8979 - 6709= 2270
#100 a=7103; b=5652; sub =1; op0=1; op1=0; // 7103 - 5652= 1451
#100 a=7992; b=8180; sub =0; op0=0; op1=1; // 7992 | 8180
#100 a=7538; b=1187; sub =0; op0=0; op1=0; // 7538 & 1187
#100 a=8827; b=2534; sub =1; op0=1; op1=0; // 8827 - 2534= 6293
#100 a=117; b=1491; sub =1; op0=1; op1=1; // 117 < 1491
#100 a=7970; b=4261; sub =0; op0=0; op1=1; // 7970 | 4261
#100 a=808; b=7373; sub =0; op0=0; op1=0; // 808 & 7373
#100 a=1492; b=3762; sub =0; op0=0; op1=1; // 1492 | 3762
#100 a=4472; b=592; sub =0; op0=0; op1=0; // 4472 & 592
#100 a=3580; b=2609; sub =0; op0=0; op1=0; // 3580 & 2609
#100 a=209; b=8367; sub =0; op0=1; op1=0; // 209 + 8367= 8576
#100 a=4380; b=4300; sub =0; op0=0; op1=1; // 4380 | 4300
#100 a=2868; b=570; sub =0; op0=1; op1=0; // 2868 + 570= 3438
#100 a=8820; b=5382; sub =1; op0=1; op1=1; // 8820 < 5382
#100 a=4243; b=7316; sub =0; op0=0; op1=1; // 4243 | 7316
#100 a=1265; b=8334; sub =0; op0=0; op1=0; // 1265 & 8334
#100 a=593; b=3662; sub =0; op0=0; op1=0; // 593 & 3662
#100 a=1669; b=7195; sub =0; op0=1; op1=0; // 1669 + 7195= 8864
#100 a=9385; b=9753; sub =0; op0=0; op1=0; // 9385 & 9753
#100 a=578; b=3136; sub =1; op0=1; op1=1; // 578 < 3136
#100 a=437; b=482; sub =0; op0=0; op1=0; // 437 & 482
#100 a=8190; b=7747; sub =0; op0=0; op1=1; // 8190 | 7747
#100 a=2104; b=1817; sub =0; op0=0; op1=0; // 2104 & 1817
#100 a=2103; b=2413; sub =0; op0=1; op1=0; // 2103 + 2413= 4516
#100 a=6443; b=311; sub =1; op0=1; op1=0; // 6443 - 311= 6132
#100 a=4478; b=3453; sub =0; op0=0; op1=0; // 4478 & 3453
#100 a=2166; b=3141; sub =1; op0=1; op1=0; // 2166 - 3141= -975
#100 a=7239; b=7353; sub =1; op0=1; op1=1; // 7239 < 7353
#100 a=4051; b=3323; sub =1; op0=1; op1=1; // 4051 < 3323
#100 a=4770; b=1583; sub =0; op0=0; op1=0; // 4770 & 1583
#100 a=7905; b=5739; sub =1; op0=1; op1=0; // 7905 - 5739= 2166
#100 a=4182; b=1258; sub =0; op0=1; op1=0; // 4182 + 1258= 5440
#100 a=7732; b=7888; sub =0; op0=0; op1=1; // 7732 | 7888
#100 a=9822; b=9172; sub =1; op0=1; op1=1; // 9822 < 9172
#100 a=9234; b=118; sub =0; op0=0; op1=1; // 9234 | 118
#100 a=8891; b=2716; sub =0; op0=1; op1=0; // 8891 + 2716= 11607
#100 a=8705; b=9132; sub =0; op0=1; op1=0; // 8705 + 9132= 17837
#100 a=285; b=6503; sub =0; op0=0; op1=1; // 285 | 6503
#100 a=1454; b=7357; sub =1; op0=1; op1=1; // 1454 < 7357
#100 a=6905; b=775; sub =0; op0=0; op1=0; // 6905 & 775
#100 a=45; b=4275; sub =0; op0=1; op1=0; // 45 + 4275= 4320
#100 a=4508; b=2641; sub =1; op0=1; op1=0; // 4508 - 2641= 1867
#100 a=444; b=3537; sub =0; op0=1; op1=0; // 444 + 3537= 3981
#100 a=9461; b=8277; sub =0; op0=0; op1=1; // 9461 | 8277
#100 a=893; b=6170; sub =0; op0=1; op1=0; // 893 + 6170= 7063
#100 a=7819; b=4934; sub =1; op0=1; op1=1; // 7819 < 4934
#100 a=5695; b=9761; sub =0; op0=0; op1=0; // 5695 & 9761
#100 a=1479; b=448; sub =0; op0=0; op1=1; // 1479 | 448
#100 a=8253; b=4291; sub =0; op0=0; op1=1; // 8253 | 4291
#100 a=5778; b=8021; sub =0; op0=0; op1=1; // 5778 | 8021
#100 a=9067; b=7596; sub =0; op0=0; op1=1; // 9067 | 7596
#100 a=3367; b=1586; sub =0; op0=1; op1=0; // 3367 + 1586= 4953
#100 a=157; b=6166; sub =0; op0=1; op1=0; // 157 + 6166= 6323
#100 a=9418; b=3426; sub =0; op0=1; op1=0; // 9418 + 3426= 12844
#100 a=1554; b=6702; sub =0; op0=0; op1=1; // 1554 | 6702
#100 a=3330; b=1897; sub =0; op0=0; op1=0; // 3330 & 1897
#100 a=8058; b=6235; sub =1; op0=1; op1=0; // 8058 - 6235= 1823
#100 a=9233; b=709; sub =1; op0=1; op1=0; // 9233 - 709= 8524
#100 a=755; b=1710; sub =1; op0=1; op1=0; // 755 - 1710= -955
#100 a=3387; b=6859; sub =0; op0=0; op1=0; // 3387 & 6859
#100 a=7872; b=3330; sub =0; op0=0; op1=1; // 7872 | 3330
#100 a=4691; b=9447; sub =0; op0=0; op1=0; // 4691 & 9447
#100 a=6738; b=7751; sub =0; op0=0; op1=1; // 6738 | 7751
#100 a=650; b=58; sub =0; op0=0; op1=1; // 650 | 58
#100 a=7967; b=2562; sub =1; op0=1; op1=0; // 7967 - 2562= 5405
#100 a=7021; b=3691; sub =0; op0=1; op1=0; // 7021 + 3691= 10712
#100 a=1101; b=1539; sub =0; op0=0; op1=1; // 1101 | 1539
#100 a=5781; b=6838; sub =1; op0=1; op1=0; // 5781 - 6838= -1057
#100 a=2847; b=8255; sub =1; op0=1; op1=1; // 2847 < 8255
#100 a=6126; b=5099; sub =1; op0=1; op1=0; // 6126 - 5099= 1027
#100 a=3730; b=237; sub =0; op0=0; op1=1; // 3730 | 237
#100 a=6586; b=1928; sub =0; op0=0; op1=1; // 6586 | 1928
#100 a=9940; b=6357; sub =0; op0=1; op1=0; // 9940 + 6357= 16297
#100 a=7279; b=9543; sub =0; op0=1; op1=0; // 7279 + 9543= 16822
#100 a=2343; b=9328; sub =0; op0=0; op1=1; // 2343 | 9328
#100 a=5241; b=4497; sub =1; op0=1; op1=0; // 5241 - 4497= 744
#100 a=7774; b=7051; sub =1; op0=1; op1=1; // 7774 < 7051
#100 a=9468; b=3468; sub =1; op0=1; op1=0; // 9468 - 3468= 6000
#100 a=7728; b=6541; sub =0; op0=1; op1=0; // 7728 + 6541= 14269
#100 a=1680; b=4042; sub =0; op0=1; op1=0; // 1680 + 4042= 5722
#100 a=5970; b=3979; sub =1; op0=1; op1=1; // 5970 < 3979
#100 a=2649; b=8820; sub =0; op0=0; op1=0; // 2649 & 8820
#100 a=8494; b=852; sub =0; op0=0; op1=0; // 8494 & 852
#100 a=9638; b=6906; sub =1; op0=1; op1=1; // 9638 < 6906
#100 a=5111; b=5694; sub =0; op0=1; op1=0; // 5111 + 5694= 10805
#100 a=9555; b=3506; sub =1; op0=1; op1=0; // 9555 - 3506= 6049
#100 a=605; b=7502; sub =0; op0=1; op1=0; // 605 + 7502= 8107
#100 a=1973; b=8073; sub =0; op0=0; op1=1; // 1973 | 8073
#100 a=8643; b=8451; sub =0; op0=0; op1=1; // 8643 | 8451
#100 a=7908; b=9261; sub =0; op0=0; op1=0; // 7908 & 9261
#100 a=6123; b=1133; sub =0; op0=0; op1=0; // 6123 & 1133
#100 a=4662; b=854; sub =0; op0=1; op1=0; // 4662 + 854= 5516
#100 a=4378; b=6446; sub =1; op0=1; op1=0; // 4378 - 6446= -2068
#100 a=3745; b=4075; sub =0; op0=1; op1=0; // 3745 + 4075= 7820
#100 a=2894; b=6678; sub =1; op0=1; op1=0; // 2894 - 6678= -3784
#100 a=7965; b=9912; sub =0; op0=0; op1=0; // 7965 & 9912
#100 a=22; b=9089; sub =1; op0=1; op1=1; // 22 < 9089
#100 a=4774; b=3703; sub =1; op0=1; op1=0; // 4774 - 3703= 1071
#100 a=3889; b=3793; sub =0; op0=0; op1=1; // 3889 | 3793
#100 a=5548; b=8893; sub =0; op0=0; op1=0; // 5548 & 8893
#100 a=3552; b=7556; sub =1; op0=1; op1=0; // 3552 - 7556= -4004
#100 a=7608; b=67; sub =0; op0=1; op1=0; // 7608 + 67= 7675
#100 a=790; b=3703; sub =0; op0=0; op1=0; // 790 & 3703
#100 a=6304; b=7874; sub =1; op0=1; op1=1; // 6304 < 7874
#100 a=4475; b=3457; sub =1; op0=1; op1=0; // 4475 - 3457= 1018
#100 a=1462; b=1680; sub =0; op0=0; op1=0; // 1462 & 1680
#100 a=6836; b=2604; sub =0; op0=0; op1=1; // 6836 | 2604
#100 a=8796; b=1288; sub =0; op0=0; op1=0; // 8796 & 1288
#100 a=7195; b=8441; sub =0; op0=1; op1=0; // 7195 + 8441= 15636
#100 a=1321; b=5280; sub =0; op0=0; op1=0; // 1321 & 5280
#100 a=4262; b=8455; sub =0; op0=1; op1=0; // 4262 + 8455= 12717
#100 a=1184; b=9978; sub =0; op0=0; op1=1; // 1184 | 9978
#100 a=5019; b=4432; sub =1; op0=1; op1=0; // 5019 - 4432= 587
#100 a=5750; b=6354; sub =0; op0=0; op1=0; // 5750 & 6354
#100 a=7175; b=8956; sub =1; op0=1; op1=1; // 7175 < 8956
#100 a=6325; b=3057; sub =0; op0=0; op1=1; // 6325 | 3057
#100 a=3920; b=3886; sub =0; op0=0; op1=0; // 3920 & 3886
#100 a=883; b=1525; sub =1; op0=1; op1=0; // 883 - 1525= -642
#100 a=7304; b=8400; sub =0; op0=0; op1=1; // 7304 | 8400
#100 a=6599; b=2; sub =0; op0=0; op1=0; // 6599 & 2
#100 a=5760; b=6496; sub =1; op0=1; op1=0; // 5760 - 6496= -736
#100 a=3444; b=4590; sub =0; op0=0; op1=1; // 3444 | 4590
#100 a=5200; b=2767; sub =1; op0=1; op1=1; // 5200 < 2767
#100 a=4066; b=2769; sub =1; op0=1; op1=0; // 4066 - 2769= 1297
#100 a=5439; b=4591; sub =1; op0=1; op1=0; // 5439 - 4591= 848
#100 a=2994; b=687; sub =0; op0=0; op1=1; // 2994 | 687
#100 a=1284; b=2653; sub =1; op0=1; op1=0; // 1284 - 2653= -1369
#100 a=122; b=155; sub =0; op0=1; op1=0; // 122 + 155= 277
#100 a=7168; b=9351; sub =0; op0=1; op1=0; // 7168 + 9351= 16519
#100 a=9438; b=6072; sub =0; op0=0; op1=1; // 9438 | 6072
#100 a=9501; b=7807; sub =1; op0=1; op1=1; // 9501 < 7807
#100 a=6393; b=4311; sub =0; op0=1; op1=0; // 6393 + 4311= 10704
#100 a=4045; b=6571; sub =1; op0=1; op1=0; // 4045 - 6571= -2526
#100 a=933; b=8416; sub =1; op0=1; op1=0; // 933 - 8416= -7483
#100 a=7914; b=5355; sub =1; op0=1; op1=1; // 7914 < 5355
#100 a=8960; b=4337; sub =1; op0=1; op1=0; // 8960 - 4337= 4623
#100 a=7265; b=9648; sub =0; op0=0; op1=0; // 7265 & 9648
#100 a=6272; b=2546; sub =0; op0=1; op1=0; // 6272 + 2546= 8818
#100 a=5128; b=6960; sub =1; op0=1; op1=1; // 5128 < 6960
#100 a=7828; b=4112; sub =0; op0=1; op1=0; // 7828 + 4112= 11940
#100 a=222; b=9128; sub =1; op0=1; op1=0; // 222 - 9128= -8906
#100 a=8329; b=7974; sub =1; op0=1; op1=0; // 8329 - 7974= 355
#100 a=3784; b=7588; sub =1; op0=1; op1=1; // 3784 < 7588
#100 a=2135; b=7989; sub =0; op0=1; op1=0; // 2135 + 7989= 10124
#100 a=3903; b=1306; sub =0; op0=1; op1=0; // 3903 + 1306= 5209
#100 a=8851; b=992; sub =0; op0=0; op1=1; // 8851 | 992
#100 a=6761; b=4997; sub =1; op0=1; op1=0; // 6761 - 4997= 1764
#100 a=840; b=1647; sub =0; op0=0; op1=1; // 840 | 1647
#100 a=9684; b=9221; sub =0; op0=0; op1=1; // 9684 | 9221
#100 a=3375; b=7983; sub =1; op0=1; op1=0; // 3375 - 7983= -4608
#100 a=7129; b=4670; sub =0; op0=1; op1=0; // 7129 + 4670= 11799
#100 a=9387; b=1537; sub =0; op0=0; op1=1; // 9387 | 1537
#100 a=7047; b=2683; sub =1; op0=1; op1=0; // 7047 - 2683= 4364
#100 a=6912; b=6476; sub =1; op0=1; op1=0; // 6912 - 6476= 436
#100 a=3341; b=7872; sub =0; op0=0; op1=0; // 3341 & 7872
#100 a=8060; b=137; sub =0; op0=1; op1=0; // 8060 + 137= 8197
#100 a=9760; b=8172; sub =0; op0=0; op1=0; // 9760 & 8172
#100 a=2745; b=7181; sub =1; op0=1; op1=1; // 2745 < 7181
#100 a=5965; b=5150; sub =1; op0=1; op1=1; // 5965 < 5150
#100 a=8754; b=4043; sub =0; op0=0; op1=1; // 8754 | 4043
#100 a=8738; b=9354; sub =0; op0=1; op1=0; // 8738 + 9354= 18092
#100 a=9189; b=4678; sub =0; op0=1; op1=0; // 9189 + 4678= 13867
#100 a=1486; b=1782; sub =0; op0=0; op1=1; // 1486 | 1782
#100 a=1795; b=8998; sub =0; op0=0; op1=1; // 1795 | 8998
#100 a=4177; b=3132; sub =1; op0=1; op1=0; // 4177 - 3132= 1045
#100 a=8515; b=8527; sub =1; op0=1; op1=1; // 8515 < 8527
#100 a=5516; b=6824; sub =1; op0=1; op1=1; // 5516 < 6824
#100 a=5018; b=4739; sub =0; op0=0; op1=0; // 5018 & 4739
#100 a=2245; b=2543; sub =0; op0=0; op1=0; // 2245 & 2543
#100 a=4067; b=7907; sub =0; op0=0; op1=0; // 4067 & 7907
#100 a=2752; b=4800; sub =0; op0=0; op1=1; // 2752 | 4800
#100 a=5102; b=8487; sub =1; op0=1; op1=0; // 5102 - 8487= -3385
#100 a=9802; b=5817; sub =0; op0=1; op1=0; // 9802 + 5817= 15619
#100 a=9075; b=8414; sub =1; op0=1; op1=0; // 9075 - 8414= 661
#100 a=2659; b=6774; sub =0; op0=0; op1=1; // 2659 | 6774
#100 a=1606; b=7470; sub =0; op0=0; op1=0; // 1606 & 7470
#100 a=4440; b=5512; sub =0; op0=0; op1=0; // 4440 & 5512
#100 a=9912; b=1106; sub =0; op0=0; op1=1; // 9912 | 1106
#100 a=1287; b=1509; sub =0; op0=0; op1=0; // 1287 & 1509
#100 a=7392; b=8521; sub =0; op0=0; op1=1; // 7392 | 8521
#100 a=2484; b=7123; sub =1; op0=1; op1=0; // 2484 - 7123= -4639
#100 a=6623; b=2819; sub =1; op0=1; op1=0; // 6623 - 2819= 3804
#100 a=1993; b=1287; sub =0; op0=0; op1=0; // 1993 & 1287
#100 a=4353; b=2539; sub =0; op0=1; op1=0; // 4353 + 2539= 6892
#100 a=9712; b=2087; sub =0; op0=0; op1=0; // 9712 & 2087
#100 a=2958; b=4887; sub =1; op0=1; op1=1; // 2958 < 4887
#100 a=7237; b=8904; sub =1; op0=1; op1=0; // 7237 - 8904= -1667
#100 a=8892; b=4781; sub =1; op0=1; op1=1; // 8892 < 4781
#100 a=8814; b=4062; sub =1; op0=1; op1=0; // 8814 - 4062= 4752
#100 a=1650; b=8179; sub =1; op0=1; op1=1; // 1650 < 8179
#100 a=6543; b=7454; sub =0; op0=0; op1=0; // 6543 & 7454
#100 a=2507; b=5039; sub =1; op0=1; op1=1; // 2507 < 5039
#100 a=4984; b=9887; sub =1; op0=1; op1=0; // 4984 - 9887= -4903
#100 a=5446; b=3698; sub =0; op0=0; op1=1; // 5446 | 3698
#100 a=4240; b=2622; sub =1; op0=1; op1=0; // 4240 - 2622= 1618
#100 a=2322; b=2129; sub =1; op0=1; op1=0; // 2322 - 2129= 193
#100 a=9953; b=5597; sub =1; op0=1; op1=0; // 9953 - 5597= 4356
#100 a=9923; b=3828; sub =1; op0=1; op1=1; // 9923 < 3828
#100 a=7902; b=2544; sub =0; op0=1; op1=0; // 7902 + 2544= 10446
#100 a=8597; b=7634; sub =1; op0=1; op1=1; // 8597 < 7634
#100 a=662; b=2200; sub =0; op0=0; op1=1; // 662 | 2200
#100 a=4575; b=7719; sub =1; op0=1; op1=1; // 4575 < 7719
#100 a=6372; b=7785; sub =0; op0=0; op1=1; // 6372 | 7785
#100 a=5863; b=139; sub =1; op0=1; op1=1; // 5863 < 139
#100 a=6412; b=7302; sub =0; op0=0; op1=1; // 6412 | 7302
#100 a=2937; b=2587; sub =0; op0=0; op1=1; // 2937 | 2587
#100 a=3135; b=3375; sub =1; op0=1; op1=1; // 3135 < 3375
#100 a=2483; b=7818; sub =0; op0=0; op1=1; // 2483 | 7818
#100 a=6984; b=5527; sub =0; op0=1; op1=0; // 6984 + 5527= 12511
#100 a=814; b=8917; sub =0; op0=0; op1=0; // 814 & 8917
#100 a=2954; b=932; sub =0; op0=0; op1=0; // 2954 & 932
#100 a=1263; b=3537; sub =1; op0=1; op1=0; // 1263 - 3537= -2274
#100 a=8874; b=4616; sub =0; op0=0; op1=0; // 8874 & 4616
#100 a=9739; b=7101; sub =0; op0=0; op1=1; // 9739 | 7101
#100 a=1754; b=8234; sub =1; op0=1; op1=0; // 1754 - 8234= -6480
#100 a=3446; b=1944; sub =1; op0=1; op1=0; // 3446 - 1944= 1502
#100 a=933; b=8474; sub =0; op0=1; op1=0; // 933 + 8474= 9407
#100 a=6731; b=8477; sub =1; op0=1; op1=0; // 6731 - 8477= -1746
#100 a=5658; b=555; sub =1; op0=1; op1=0; // 5658 - 555= 5103
#100 a=3431; b=1780; sub =0; op0=1; op1=0; // 3431 + 1780= 5211
#100 a=7944; b=3265; sub =0; op0=0; op1=0; // 7944 & 3265
#100 a=3819; b=9319; sub =0; op0=1; op1=0; // 3819 + 9319= 13138
#100 a=4425; b=1869; sub =1; op0=1; op1=1; // 4425 < 1869
#100 a=9402; b=5286; sub =0; op0=0; op1=0; // 9402 & 5286
#100 a=3285; b=5026; sub =1; op0=1; op1=1; // 3285 < 5026
#100 a=8170; b=3182; sub =0; op0=0; op1=0; // 8170 & 3182
#100 a=347; b=8974; sub =0; op0=1; op1=0; // 347 + 8974= 9321
#100 a=2698; b=4586; sub =1; op0=1; op1=1; // 2698 < 4586
#100 a=7382; b=8319; sub =0; op0=0; op1=1; // 7382 | 8319
#100 a=1896; b=7479; sub =1; op0=1; op1=0; // 1896 - 7479= -5583
#100 a=7563; b=6672; sub =1; op0=1; op1=0; // 7563 - 6672= 891
#100 a=2146; b=2307; sub =0; op0=0; op1=1; // 2146 | 2307
#100 a=6147; b=9063; sub =1; op0=1; op1=0; // 6147 - 9063= -2916
#100 a=9616; b=2944; sub =0; op0=0; op1=0; // 9616 & 2944
#100 a=1278; b=9700; sub =1; op0=1; op1=1; // 1278 < 9700
#100 a=3803; b=4160; sub =1; op0=1; op1=0; // 3803 - 4160= -357
#100 a=9407; b=291; sub =0; op0=0; op1=0; // 9407 & 291
#100 a=3188; b=1641; sub =0; op0=0; op1=1; // 3188 | 1641
#100 a=9987; b=4593; sub =1; op0=1; op1=1; // 9987 < 4593
#100 a=164; b=4491; sub =0; op0=0; op1=1; // 164 | 4491
#100 a=9668; b=9939; sub =1; op0=1; op1=0; // 9668 - 9939= -271
#100 a=6593; b=7859; sub =0; op0=0; op1=1; // 6593 | 7859
#100 a=7690; b=43; sub =1; op0=1; op1=0; // 7690 - 43= 7647
#100 a=424; b=7297; sub =0; op0=0; op1=0; // 424 & 7297
#100 a=9168; b=766; sub =0; op0=1; op1=0; // 9168 + 766= 9934
#100 a=3459; b=3568; sub =0; op0=0; op1=0; // 3459 & 3568
#100 a=2381; b=3051; sub =0; op0=1; op1=0; // 2381 + 3051= 5432
#100 a=5879; b=2208; sub =1; op0=1; op1=0; // 5879 - 2208= 3671
#100 a=2895; b=3775; sub =0; op0=0; op1=0; // 2895 & 3775
#100 a=8232; b=4042; sub =1; op0=1; op1=1; // 8232 < 4042
#100 a=65; b=781; sub =1; op0=1; op1=0; // 65 - 781= -716
#100 a=8005; b=9957; sub =1; op0=1; op1=1; // 8005 < 9957
#100 a=7766; b=3141; sub =1; op0=1; op1=0; // 7766 - 3141= 4625
#100 a=6093; b=3415; sub =0; op0=0; op1=1; // 6093 | 3415
#100 a=3305; b=6727; sub =0; op0=0; op1=1; // 3305 | 6727
#100 a=4190; b=9251; sub =0; op0=0; op1=1; // 4190 | 9251
#100 a=4585; b=388; sub =0; op0=0; op1=1; // 4585 | 388
#100 a=8739; b=7197; sub =0; op0=0; op1=0; // 8739 & 7197
#100 a=239; b=2756; sub =0; op0=0; op1=0; // 239 & 2756
#100 a=9790; b=7765; sub =0; op0=0; op1=0; // 9790 & 7765
#100 a=5413; b=8610; sub =0; op0=0; op1=0; // 5413 & 8610
#100 a=3723; b=5884; sub =1; op0=1; op1=1; // 3723 < 5884
#100 a=2498; b=1625; sub =0; op0=0; op1=1; // 2498 | 1625
#100 a=3060; b=9098; sub =1; op0=1; op1=0; // 3060 - 9098= -6038
#100 a=3575; b=9286; sub =1; op0=1; op1=1; // 3575 < 9286
#100 a=9685; b=99; sub =1; op0=1; op1=1; // 9685 < 99
#100 a=8816; b=3487; sub =0; op0=0; op1=1; // 8816 | 3487
#100 a=3759; b=4623; sub =0; op0=0; op1=0; // 3759 & 4623
#100 a=9984; b=7137; sub =1; op0=1; op1=1; // 9984 < 7137
#100 a=1790; b=3356; sub =1; op0=1; op1=1; // 1790 < 3356
#100 a=9721; b=2636; sub =0; op0=0; op1=0; // 9721 & 2636
#100 a=3563; b=1497; sub =0; op0=1; op1=0; // 3563 + 1497= 5060
#100 a=19; b=1637; sub =0; op0=0; op1=1; // 19 | 1637
#100 a=2949; b=3784; sub =0; op0=0; op1=0; // 2949 & 3784
#100 a=6373; b=8353; sub =0; op0=0; op1=1; // 6373 | 8353
#100 a=8617; b=8148; sub =0; op0=0; op1=0; // 8617 & 8148
#100 a=1541; b=6539; sub =1; op0=1; op1=1; // 1541 < 6539
#100 a=447; b=5602; sub =1; op0=1; op1=0; // 447 - 5602= -5155
#100 a=4405; b=1763; sub =1; op0=1; op1=0; // 4405 - 1763= 2642
#100 a=1919; b=6356; sub =1; op0=1; op1=1; // 1919 < 6356
#100 a=7779; b=1462; sub =0; op0=0; op1=1; // 7779 | 1462
#100 a=2581; b=1990; sub =1; op0=1; op1=1; // 2581 < 1990
#100 a=1445; b=1090; sub =1; op0=1; op1=0; // 1445 - 1090= 355
#100 a=6811; b=3429; sub =1; op0=1; op1=1; // 6811 < 3429
#100 a=1582; b=3070; sub =0; op0=0; op1=1; // 1582 | 3070
#100 a=2690; b=1886; sub =1; op0=1; op1=0; // 2690 - 1886= 804
#100 a=1238; b=8808; sub =1; op0=1; op1=0; // 1238 - 8808= -7570
#100 a=7981; b=9091; sub =1; op0=1; op1=1; // 7981 < 9091
#100 a=4401; b=4541; sub =0; op0=1; op1=0; // 4401 + 4541= 8942
#100 a=1533; b=5217; sub =0; op0=0; op1=0; // 1533 & 5217
#100 a=6737; b=2477; sub =1; op0=1; op1=0; // 6737 - 2477= 4260
#100 a=8957; b=4651; sub =1; op0=1; op1=0; // 8957 - 4651= 4306
#100 a=2552; b=4008; sub =1; op0=1; op1=1; // 2552 < 4008
#100 a=4414; b=2869; sub =0; op0=1; op1=0; // 4414 + 2869= 7283
#100 a=9225; b=4107; sub =1; op0=1; op1=1; // 9225 < 4107
#100 a=1579; b=8062; sub =0; op0=1; op1=0; // 1579 + 8062= 9641
#100 a=7570; b=2371; sub =0; op0=1; op1=0; // 7570 + 2371= 9941
#100 a=3110; b=2595; sub =1; op0=1; op1=0; // 3110 - 2595= 515
#100 a=1209; b=6448; sub =1; op0=1; op1=0; // 1209 - 6448= -5239
#100 a=1081; b=9249; sub =0; op0=1; op1=0; // 1081 + 9249= 10330
#100 a=6735; b=7996; sub =0; op0=1; op1=0; // 6735 + 7996= 14731
#100 a=7617; b=1075; sub =1; op0=1; op1=1; // 7617 < 1075
#100 a=747; b=7920; sub =0; op0=0; op1=1; // 747 | 7920
#100 a=3977; b=9955; sub =0; op0=0; op1=1; // 3977 | 9955
#100 a=3846; b=1182; sub =0; op0=0; op1=0; // 3846 & 1182
#100 a=2217; b=2177; sub =0; op0=0; op1=0; // 2217 & 2177
#100 a=3831; b=4694; sub =0; op0=1; op1=0; // 3831 + 4694= 8525
#100 a=2486; b=285; sub =0; op0=0; op1=0; // 2486 & 285
#100 a=7830; b=2713; sub =0; op0=1; op1=0; // 7830 + 2713= 10543
#100 a=6057; b=8933; sub =0; op0=0; op1=1; // 6057 | 8933
#100 a=6646; b=9093; sub =0; op0=1; op1=0; // 6646 + 9093= 15739
#100 a=9252; b=903; sub =1; op0=1; op1=1; // 9252 < 903
#100 a=9701; b=9259; sub =1; op0=1; op1=1; // 9701 < 9259
#100 a=9296; b=6288; sub =1; op0=1; op1=1; // 9296 < 6288
#100 a=7335; b=1227; sub =0; op0=1; op1=0; // 7335 + 1227= 8562
#100 a=6823; b=791; sub =0; op0=1; op1=0; // 6823 + 791= 7614
#100 a=5491; b=6457; sub =0; op0=0; op1=0; // 5491 & 6457
#100 a=10; b=3788; sub =0; op0=0; op1=1; // 10 | 3788
#100 a=1748; b=9774; sub =1; op0=1; op1=0; // 1748 - 9774= -8026
#100 a=4114; b=154; sub =0; op0=0; op1=0; // 4114 & 154
#100 a=3946; b=5602; sub =0; op0=0; op1=1; // 3946 | 5602
#100 a=8532; b=8468; sub =0; op0=0; op1=1; // 8532 | 8468
#100 a=1450; b=7749; sub =1; op0=1; op1=0; // 1450 - 7749= -6299
#100 a=4374; b=1046; sub =0; op0=0; op1=0; // 4374 & 1046
#100 a=2472; b=2174; sub =1; op0=1; op1=0; // 2472 - 2174= 298
#100 a=6897; b=6129; sub =1; op0=1; op1=0; // 6897 - 6129= 768
#100 a=3311; b=5160; sub =0; op0=0; op1=1; // 3311 | 5160
#100 a=7020; b=5326; sub =0; op0=0; op1=0; // 7020 & 5326
#100 a=7545; b=3857; sub =0; op0=1; op1=0; // 7545 + 3857= 11402
#100 a=1875; b=3770; sub =1; op0=1; op1=0; // 1875 - 3770= -1895
#100 a=771; b=3016; sub =0; op0=0; op1=0; // 771 & 3016
#100 a=7467; b=7765; sub =1; op0=1; op1=0; // 7467 - 7765= -298
#100 a=1262; b=5512; sub =0; op0=0; op1=0; // 1262 & 5512
#100 a=8565; b=7799; sub =0; op0=1; op1=0; // 8565 + 7799= 16364
#100 a=7859; b=2480; sub =0; op0=0; op1=1; // 7859 | 2480
#100 a=9248; b=8881; sub =0; op0=0; op1=0; // 9248 & 8881
#100 a=1907; b=6606; sub =0; op0=0; op1=0; // 1907 & 6606
#100 a=6714; b=8171; sub =0; op0=0; op1=1; // 6714 | 8171
#100 a=8277; b=1690; sub =0; op0=1; op1=0; // 8277 + 1690= 9967
#100 a=6848; b=8749; sub =1; op0=1; op1=0; // 6848 - 8749= -1901
#100 a=6143; b=7522; sub =0; op0=0; op1=1; // 6143 | 7522
#100 a=5946; b=2530; sub =0; op0=0; op1=0; // 5946 & 2530
#100 a=7881; b=3060; sub =0; op0=1; op1=0; // 7881 + 3060= 10941
#100 a=7741; b=5867; sub =0; op0=0; op1=1; // 7741 | 5867
#100 a=3761; b=6906; sub =0; op0=0; op1=1; // 3761 | 6906
#100 a=1901; b=1385; sub =1; op0=1; op1=1; // 1901 < 1385
#100 a=932; b=4739; sub =1; op0=1; op1=1; // 932 < 4739
#100 a=805; b=9833; sub =1; op0=1; op1=0; // 805 - 9833= -9028
#100 a=4548; b=2016; sub =0; op0=0; op1=1; // 4548 | 2016
#100 a=7016; b=8844; sub =0; op0=1; op1=0; // 7016 + 8844= 15860
#100 a=5299; b=5172; sub =0; op0=1; op1=0; // 5299 + 5172= 10471
#100 a=9547; b=4393; sub =0; op0=0; op1=0; // 9547 & 4393
#100 a=6592; b=6550; sub =0; op0=1; op1=0; // 6592 + 6550= 13142
#100 a=256; b=3499; sub =1; op0=1; op1=0; // 256 - 3499= -3243
#100 a=9118; b=4136; sub =0; op0=0; op1=1; // 9118 | 4136
#100 a=1799; b=1874; sub =0; op0=0; op1=0; // 1799 & 1874
#100 a=8199; b=6499; sub =1; op0=1; op1=1; // 8199 < 6499
#100 a=1616; b=3777; sub =0; op0=1; op1=0; // 1616 + 3777= 5393
#100 a=9806; b=364; sub =0; op0=0; op1=1; // 9806 | 364
#100 a=5262; b=7698; sub =0; op0=0; op1=1; // 5262 | 7698
#100 a=9371; b=5765; sub =1; op0=1; op1=1; // 9371 < 5765
#100 a=4452; b=1153; sub =0; op0=1; op1=0; // 4452 + 1153= 5605
#100 a=2296; b=8777; sub =1; op0=1; op1=0; // 2296 - 8777= -6481
#100 a=7494; b=5160; sub =0; op0=0; op1=1; // 7494 | 5160
#100 a=1209; b=1514; sub =0; op0=0; op1=0; // 1209 & 1514
#100 a=3829; b=9681; sub =1; op0=1; op1=1; // 3829 < 9681
#100 a=3538; b=3794; sub =1; op0=1; op1=0; // 3538 - 3794= -256
#100 a=1663; b=4254; sub =1; op0=1; op1=1; // 1663 < 4254
#100 a=6644; b=6145; sub =0; op0=0; op1=0; // 6644 & 6145
#100 a=3254; b=9048; sub =0; op0=0; op1=1; // 3254 | 9048
#100 a=4710; b=5926; sub =0; op0=0; op1=0; // 4710 & 5926
#100 a=6925; b=2547; sub =0; op0=0; op1=1; // 6925 | 2547
#100 a=7567; b=4596; sub =0; op0=0; op1=0; // 7567 & 4596
#100 a=3113; b=8319; sub =1; op0=1; op1=1; // 3113 < 8319
#100 a=7946; b=7497; sub =0; op0=1; op1=0; // 7946 + 7497= 15443
#100 a=4978; b=4584; sub =1; op0=1; op1=0; // 4978 - 4584= 394
#100 a=5751; b=5955; sub =1; op0=1; op1=0; // 5751 - 5955= -204
#100 a=6158; b=534; sub =0; op0=0; op1=1; // 6158 | 534
#100 a=4991; b=3208; sub =0; op0=1; op1=0; // 4991 + 3208= 8199
#100 a=5728; b=2963; sub =0; op0=1; op1=0; // 5728 + 2963= 8691
#100 a=8768; b=314; sub =0; op0=1; op1=0; // 8768 + 314= 9082
#100 a=877; b=8523; sub =0; op0=0; op1=1; // 877 | 8523
#100 a=7777; b=5937; sub =0; op0=0; op1=0; // 7777 & 5937
#100 a=4551; b=9655; sub =0; op0=0; op1=0; // 4551 & 9655
#100 a=7213; b=5118; sub =1; op0=1; op1=0; // 7213 - 5118= 2095
#100 a=1656; b=4180; sub =1; op0=1; op1=0; // 1656 - 4180= -2524
#100 a=5313; b=4175; sub =1; op0=1; op1=0; // 5313 - 4175= 1138
#100 a=7175; b=1004; sub =1; op0=1; op1=0; // 7175 - 1004= 6171
#100 a=6563; b=9441; sub =1; op0=1; op1=0; // 6563 - 9441= -2878
#100 a=6654; b=9978; sub =0; op0=0; op1=1; // 6654 | 9978
#100 a=6042; b=1338; sub =1; op0=1; op1=0; // 6042 - 1338= 4704
#100 a=7622; b=7372; sub =0; op0=0; op1=1; // 7622 | 7372
#100 a=1713; b=9637; sub =0; op0=0; op1=1; // 1713 | 9637
#100 a=1004; b=4962; sub =0; op0=0; op1=0; // 1004 & 4962
#100 a=434; b=4703; sub =1; op0=1; op1=1; // 434 < 4703
#100 a=5248; b=5371; sub =0; op0=1; op1=0; // 5248 + 5371= 10619
#100 a=8449; b=7368; sub =1; op0=1; op1=1; // 8449 < 7368
#100 a=147; b=757; sub =0; op0=0; op1=0; // 147 & 757
#100 a=6264; b=1237; sub =0; op0=0; op1=0; // 6264 & 1237
#100 a=7927; b=5899; sub =0; op0=1; op1=0; // 7927 + 5899= 13826
#100 a=4643; b=6798; sub =0; op0=0; op1=1; // 4643 | 6798
#100 a=4974; b=2835; sub =0; op0=0; op1=1; // 4974 | 2835
#100 a=6685; b=9299; sub =0; op0=0; op1=1; // 6685 | 9299
#100 a=3371; b=2167; sub =1; op0=1; op1=1; // 3371 < 2167
#100 a=1614; b=9764; sub =0; op0=0; op1=1; // 1614 | 9764
#100 a=3355; b=8465; sub =0; op0=0; op1=1; // 3355 | 8465
#100 a=7694; b=5699; sub =0; op0=0; op1=1; // 7694 | 5699
#100 a=8361; b=6069; sub =1; op0=1; op1=1; // 8361 < 6069
#100 a=1103; b=7423; sub =0; op0=0; op1=0; // 1103 & 7423
#100 a=6017; b=3514; sub =1; op0=1; op1=1; // 6017 < 3514
#100 a=2956; b=4190; sub =1; op0=1; op1=1; // 2956 < 4190
#100 a=601; b=2461; sub =0; op0=1; op1=0; // 601 + 2461= 3062
#100 a=2338; b=6022; sub =0; op0=0; op1=0; // 2338 & 6022
#100 a=6820; b=3166; sub =0; op0=1; op1=0; // 6820 + 3166= 9986
#100 a=8154; b=9201; sub =0; op0=0; op1=0; // 8154 & 9201
#100 a=5047; b=8484; sub =0; op0=0; op1=1; // 5047 | 8484
#100 a=2532; b=7888; sub =0; op0=1; op1=0; // 2532 + 7888= 10420
#100 a=722; b=4985; sub =0; op0=0; op1=1; // 722 | 4985
#100 a=1744; b=4; sub =0; op0=0; op1=1; // 1744 | 4
#100 a=2494; b=6746; sub =0; op0=1; op1=0; // 2494 + 6746= 9240
#100 a=3484; b=1442; sub =1; op0=1; op1=0; // 3484 - 1442= 2042
#100 a=9994; b=3752; sub =0; op0=0; op1=0; // 9994 & 3752
#100 a=8504; b=5730; sub =1; op0=1; op1=0; // 8504 - 5730= 2774
#100 a=7542; b=236; sub =0; op0=0; op1=1; // 7542 | 236
#100 a=5798; b=7876; sub =0; op0=0; op1=0; // 5798 & 7876
#100 a=1253; b=667; sub =0; op0=1; op1=0; // 1253 + 667= 1920
#100 a=9353; b=9429; sub =0; op0=0; op1=1; // 9353 | 9429
#100 a=603; b=6631; sub =0; op0=0; op1=0; // 603 & 6631
#100 a=1706; b=5382; sub =0; op0=1; op1=0; // 1706 + 5382= 7088
#100 a=406; b=5023; sub =1; op0=1; op1=0; // 406 - 5023= -4617
#100 a=324; b=8301; sub =0; op0=0; op1=1; // 324 | 8301
#100 a=2999; b=5159; sub =0; op0=0; op1=0; // 2999 & 5159
#100 a=8226; b=1913; sub =0; op0=0; op1=1; // 8226 | 1913
#100 a=4122; b=8700; sub =0; op0=0; op1=1; // 4122 | 8700
#100 a=964; b=3406; sub =0; op0=0; op1=0; // 964 & 3406
#100 a=3896; b=5824; sub =1; op0=1; op1=0; // 3896 - 5824= -1928
#100 a=4563; b=2910; sub =0; op0=0; op1=1; // 4563 | 2910
#100 a=61; b=6076; sub =0; op0=1; op1=0; // 61 + 6076= 6137
#100 a=8396; b=2666; sub =1; op0=1; op1=1; // 8396 < 2666
#100 a=4130; b=185; sub =1; op0=1; op1=1; // 4130 < 185
#100 a=628; b=2216; sub =0; op0=1; op1=0; // 628 + 2216= 2844
#100 a=8618; b=7406; sub =1; op0=1; op1=1; // 8618 < 7406
#100 a=5752; b=843; sub =0; op0=0; op1=1; // 5752 | 843
#100 a=4234; b=834; sub =1; op0=1; op1=0; // 4234 - 834= 3400
#100 a=2928; b=4082; sub =0; op0=0; op1=1; // 2928 | 4082
#100 a=9850; b=1252; sub =0; op0=1; op1=0; // 9850 + 1252= 11102
#100 a=4722; b=3290; sub =0; op0=0; op1=1; // 4722 | 3290
#100 a=6737; b=2126; sub =1; op0=1; op1=0; // 6737 - 2126= 4611
#100 a=1528; b=881; sub =1; op0=1; op1=1; // 1528 < 881
#100 a=2365; b=674; sub =1; op0=1; op1=1; // 2365 < 674
#100 a=799; b=4689; sub =0; op0=0; op1=0; // 799 & 4689
#100 a=3495; b=7976; sub =0; op0=1; op1=0; // 3495 + 7976= 11471
#100 a=3677; b=3442; sub =0; op0=0; op1=1; // 3677 | 3442
#100 a=500; b=5237; sub =0; op0=1; op1=0; // 500 + 5237= 5737
#100 a=9883; b=5089; sub =1; op0=1; op1=0; // 9883 - 5089= 4794
#100 a=4861; b=7807; sub =0; op0=1; op1=0; // 4861 + 7807= 12668
#100 a=4904; b=2707; sub =0; op0=1; op1=0; // 4904 + 2707= 7611
#100 a=5232; b=9195; sub =0; op0=0; op1=1; // 5232 | 9195
#100 a=9677; b=4461; sub =1; op0=1; op1=0; // 9677 - 4461= 5216
#100 a=6809; b=8999; sub =0; op0=0; op1=1; // 6809 | 8999
#100 a=2962; b=8700; sub =1; op0=1; op1=0; // 2962 - 8700= -5738
#100 a=6425; b=2748; sub =0; op0=0; op1=0; // 6425 & 2748
#100 a=878; b=3577; sub =0; op0=0; op1=0; // 878 & 3577
#100 a=5065; b=6965; sub =0; op0=1; op1=0; // 5065 + 6965= 12030
#100 a=3411; b=7881; sub =0; op0=0; op1=0; // 3411 & 7881
#100 a=658; b=8128; sub =0; op0=0; op1=0; // 658 & 8128
#100 a=6528; b=9775; sub =1; op0=1; op1=0; // 6528 - 9775= -3247
#100 a=2615; b=3011; sub =0; op0=0; op1=1; // 2615 | 3011
#100 a=4597; b=6654; sub =1; op0=1; op1=0; // 4597 - 6654= -2057
#100 a=3910; b=2695; sub =0; op0=0; op1=1; // 3910 | 2695
#100 a=4253; b=2573; sub =0; op0=0; op1=0; // 4253 & 2573
#100 a=7051; b=2469; sub =1; op0=1; op1=0; // 7051 - 2469= 4582
#100 a=4143; b=5210; sub =1; op0=1; op1=1; // 4143 < 5210
#100 a=1537; b=8942; sub =0; op0=1; op1=0; // 1537 + 8942= 10479
#100 a=333; b=8589; sub =1; op0=1; op1=0; // 333 - 8589= -8256
#100 a=2790; b=6542; sub =0; op0=0; op1=1; // 2790 | 6542
#100 a=1551; b=7801; sub =1; op0=1; op1=1; // 1551 < 7801
#100 a=3376; b=389; sub =0; op0=0; op1=1; // 3376 | 389
#100 a=717; b=9910; sub =0; op0=0; op1=0; // 717 & 9910
#100 a=336; b=5380; sub =1; op0=1; op1=1; // 336 < 5380
#100 a=3908; b=8922; sub =1; op0=1; op1=0; // 3908 - 8922= -5014
#100 a=6945; b=973; sub =0; op0=0; op1=1; // 6945 | 973
#100 a=4853; b=3784; sub =0; op0=1; op1=0; // 4853 + 3784= 8637
#100 a=9385; b=1049; sub =0; op0=1; op1=0; // 9385 + 1049= 10434
#100 a=9799; b=8680; sub =0; op0=1; op1=0; // 9799 + 8680= 18479
#100 a=1497; b=4537; sub =0; op0=0; op1=0; // 1497 & 4537
#100 a=6120; b=5605; sub =0; op0=1; op1=0; // 6120 + 5605= 11725
#100 a=8918; b=9417; sub =1; op0=1; op1=1; // 8918 < 9417
#100 a=5984; b=8125; sub =0; op0=1; op1=0; // 5984 + 8125= 14109
#100 a=6510; b=6384; sub =0; op0=1; op1=0; // 6510 + 6384= 12894
#100 a=3634; b=7955; sub =0; op0=1; op1=0; // 3634 + 7955= 11589
#100 a=7232; b=423; sub =0; op0=0; op1=1; // 7232 | 423
#100 a=3602; b=2895; sub =0; op0=1; op1=0; // 3602 + 2895= 6497
#100 a=533; b=5481; sub =0; op0=1; op1=0; // 533 + 5481= 6014
#100 a=651; b=2707; sub =1; op0=1; op1=0; // 651 - 2707= -2056
#100 a=6837; b=4230; sub =1; op0=1; op1=1; // 6837 < 4230
#100 a=5586; b=8209; sub =1; op0=1; op1=1; // 5586 < 8209
#100 a=6590; b=6979; sub =1; op0=1; op1=0; // 6590 - 6979= -389
#100 a=5918; b=8949; sub =0; op0=0; op1=0; // 5918 & 8949
#100 a=9093; b=976; sub =0; op0=0; op1=0; // 9093 & 976
#100 a=148; b=6178; sub =1; op0=1; op1=1; // 148 < 6178
#100 a=3182; b=9959; sub =1; op0=1; op1=0; // 3182 - 9959= -6777
#100 a=5772; b=2947; sub =1; op0=1; op1=0; // 5772 - 2947= 2825
#100 a=474; b=9454; sub =1; op0=1; op1=1; // 474 < 9454
#100 a=663; b=9662; sub =0; op0=0; op1=1; // 663 | 9662
#100 a=2689; b=9594; sub =0; op0=1; op1=0; // 2689 + 9594= 12283
#100 a=5741; b=9646; sub =0; op0=0; op1=1; // 5741 | 9646
#100 a=6160; b=2007; sub =0; op0=1; op1=0; // 6160 + 2007= 8167
#100 a=7363; b=7715; sub =0; op0=1; op1=0; // 7363 + 7715= 15078
#100 a=4296; b=6675; sub =0; op0=1; op1=0; // 4296 + 6675= 10971
#100 a=5534; b=7798; sub =0; op0=0; op1=0; // 5534 & 7798
#100 a=7117; b=8241; sub =0; op0=1; op1=0; // 7117 + 8241= 15358
#100 a=9039; b=9439; sub =0; op0=1; op1=0; // 9039 + 9439= 18478
#100 a=3724; b=5699; sub =0; op0=0; op1=1; // 3724 | 5699
#100 a=9108; b=7325; sub =0; op0=1; op1=0; // 9108 + 7325= 16433
#100 a=7500; b=8285; sub =1; op0=1; op1=0; // 7500 - 8285= -785
#100 a=8244; b=3641; sub =0; op0=1; op1=0; // 8244 + 3641= 11885
#100 a=2663; b=6238; sub =0; op0=0; op1=1; // 2663 | 6238
#100 a=5197; b=6515; sub =0; op0=1; op1=0; // 5197 + 6515= 11712
#100 a=1767; b=210; sub =1; op0=1; op1=0; // 1767 - 210= 1557
#100 a=6467; b=2655; sub =0; op0=0; op1=0; // 6467 & 2655
#100 a=4769; b=8094; sub =1; op0=1; op1=1; // 4769 < 8094
#100 a=3447; b=8727; sub =1; op0=1; op1=0; // 3447 - 8727= -5280
#100 a=9233; b=2852; sub =1; op0=1; op1=0; // 9233 - 2852= 6381
#100 a=4130; b=5270; sub =1; op0=1; op1=0; // 4130 - 5270= -1140
#100 a=6903; b=7219; sub =0; op0=1; op1=0; // 6903 + 7219= 14122
#100 a=1310; b=9282; sub =0; op0=0; op1=0; // 1310 & 9282
#100 a=8326; b=1145; sub =1; op0=1; op1=0; // 8326 - 1145= 7181
#100 a=7410; b=9065; sub =1; op0=1; op1=1; // 7410 < 9065
#100 a=1464; b=6375; sub =0; op0=0; op1=0; // 1464 & 6375
#100 a=2179; b=3898; sub =0; op0=0; op1=0; // 2179 & 3898
#100 a=9367; b=8262; sub =1; op0=1; op1=0; // 9367 - 8262= 1105
#100 a=2285; b=684; sub =0; op0=0; op1=0; // 2285 & 684
#100 a=6770; b=1995; sub =1; op0=1; op1=1; // 6770 < 1995
#100 a=173; b=854; sub =0; op0=1; op1=0; // 173 + 854= 1027
#100 a=4813; b=595; sub =0; op0=0; op1=1; // 4813 | 595
#100 a=4726; b=3718; sub =1; op0=1; op1=1; // 4726 < 3718
#100 a=386; b=2273; sub =0; op0=0; op1=0; // 386 & 2273
#100 a=1643; b=3459; sub =1; op0=1; op1=1; // 1643 < 3459
#100 a=4458; b=1064; sub =1; op0=1; op1=1; // 4458 < 1064
#100 a=169; b=9360; sub =0; op0=1; op1=0; // 169 + 9360= 9529
#100 a=852; b=5746; sub =0; op0=1; op1=0; // 852 + 5746= 6598
#100 a=9202; b=6299; sub =0; op0=0; op1=1; // 9202 | 6299
#100 a=5507; b=710; sub =1; op0=1; op1=0; // 5507 - 710= 4797
#100 a=2292; b=4411; sub =0; op0=0; op1=1; // 2292 | 4411
#100 a=518; b=2551; sub =1; op0=1; op1=0; // 518 - 2551= -2033
#100 a=1326; b=9487; sub =1; op0=1; op1=1; // 1326 < 9487
#100 a=2462; b=272; sub =0; op0=0; op1=1; // 2462 | 272
#100 a=2788; b=5819; sub =0; op0=0; op1=0; // 2788 & 5819
#100 a=2397; b=5408; sub =0; op0=1; op1=0; // 2397 + 5408= 7805
#100 a=5992; b=8690; sub =0; op0=0; op1=1; // 5992 | 8690
#100 a=9012; b=4446; sub =1; op0=1; op1=1; // 9012 < 4446
#100 a=6946; b=205; sub =0; op0=0; op1=0; // 6946 & 205
#100 a=7140; b=4218; sub =1; op0=1; op1=0; // 7140 - 4218= 2922


  
 #100 // Required for iverilog to show final values
 $display($time,,,, "a=%b, b=%b, sub=%b, op0=%b, op1=%b, out=%b",a,b,sub,op0,op1,out);
 end
endmodule 